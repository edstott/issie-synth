

    module RAM1_249(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 2024;
ram[1] = 35857;
ram[2] = 39169;
ram[3] = 47113;
ram[4] = 49850;
ram[5] = 63010;
ram[6] = 24584;
ram[7] = 16395;
ram[8] = 20492;
ram[9] = 16395;
ram[10] = 4660;
ram[11] = 28672;
ram[12] = 5153;
ram[13] = 28672;
ram[292] = 564;
ram[2730] = 205;
ram[2731] = 171;
ram[2733] = 17;
    end
    endmodule

    
module main (
	clk,
	RAMOUT_262_out0,
	IROUT_350_out0,
	R0OUT_38_out0,
	R1OUT_49_out0,
	R3OUT_127_out0,
	R2OUT_163_out0,
	STALL0_352_out0,
	STALLF_182_out0,
	FETCH_569_out0);
input clk;
output  [15:0] IROUT_350_out0;
output  [15:0] R0OUT_38_out0;
output  [15:0] R1OUT_49_out0;
output  [15:0] R2OUT_163_out0;
output  [15:0] R3OUT_127_out0;
output  [15:0] RAMOUT_262_out0;
output FETCH_569_out0;
output STALL0_352_out0;
output STALLF_182_out0;
reg  [11:0] REG1_274_out0 = 12'h0;
reg  [15:0] REG0_543_out0 = 16'h0;
reg  [15:0] REG1_164_out0 = 16'h0;
reg  [15:0] REG1_50_out0 = 16'h0;
reg  [15:0] REG1_51_out0 = 16'h0;
reg  [15:0] REG2_584_out0 = 16'h0;
reg  [15:0] REG3_333_out0 = 16'h0;
reg  [1:0] REG1_156_out0 = 2'h0;
reg FF1_251_out0 = 1'b0;
reg FF1_459_out0 = 1'b0;
reg FF1_538_out0 = 1'b0;
reg FF2_128_out0 = 1'b0;
reg FF2_621_out0 = 1'b0;
reg N_564_out0 = 1'b0;
reg Z_361_out0 = 1'b0;
wire  [10:0] C1_367_out0;
wire  [10:0] v_58_out0;
wire  [10:0] v_79_out0;
wire  [11:0] A1_225_out0;
wire  [11:0] A1_407_out0;
wire  [11:0] A1_8_out0;
wire  [11:0] C2_550_out0;
wire  [11:0] C2_579_out0;
wire  [11:0] C3_431_out0;
wire  [11:0] IN14_450_out0;
wire  [11:0] IN1_465_out0;
wire  [11:0] MUX1_272_out0;
wire  [11:0] MUX1_392_out0;
wire  [11:0] MUX2_642_out0;
wire  [11:0] MUX3_205_out0;
wire  [11:0] MUX5_458_out0;
wire  [11:0] MUX6_69_out0;
wire  [11:0] N_456_out0;
wire  [11:0] N_587_out0;
wire  [11:0] PCOUT_637_out0;
wire  [11:0] RAMADDRMUX_160_out0;
wire  [11:0] RAMADDRMUX_20_out0;
wire  [11:0] XOR1_588_out0;
wire  [11:0] v_102_out0;
wire  [11:0] v_285_out0;
wire  [11:0] v_320_out0;
wire  [11:0] v_489_out1;
wire  [11:0] v_499_out0;
wire  [11:0] v_623_out0;
wire  [11:0] v_74_out0;
wire  [11:0] v_89_out0;
wire  [12:0] v_319_out0;
wire  [12:0] v_412_out0;
wire  [13:0] IN14_189_out0;
wire  [13:0] IN1_257_out0;
wire  [13:0] v_145_out0;
wire  [13:0] v_25_out0;
wire  [13:0] v_339_out1;
wire  [13:0] v_566_out0;
wire  [14:0] IN14_442_out0;
wire  [14:0] IN14_610_out0;
wire  [14:0] IN1_41_out0;
wire  [14:0] IN1_477_out0;
wire  [14:0] v_151_out0;
wire  [14:0] v_18_out0;
wire  [14:0] v_293_out1;
wire  [14:0] v_42_out0;
wire  [14:0] v_48_out0;
wire  [14:0] v_52_out0;
wire  [15:0] A1_597_out0;
wire  [15:0] ALUOUT_240_out0;
wire  [15:0] ALUOUT_401_out0;
wire  [15:0] ALUOUT_503_out0;
wire  [15:0] ALUOUT_554_out0;
wire  [15:0] A_366_out0;
wire  [15:0] A_493_out0;
wire  [15:0] A_568_out0;
wire  [15:0] A_65_out0;
wire  [15:0] B_464_out0;
wire  [15:0] C1_544_out0;
wire  [15:0] DIN3_461_out0;
wire  [15:0] DIN_173_out0;
wire  [15:0] DIN_203_out0;
wire  [15:0] DIN_204_out0;
wire  [15:0] DM1_510_out0;
wire  [15:0] DM1_510_out1;
wire  [15:0] DOUT1_107_out0;
wire  [15:0] DOUT2_118_out0;
wire  [15:0] DOUT_138_out0;
wire  [15:0] DOUT_139_out0;
wire  [15:0] IN_143_out0;
wire  [15:0] IN_358_out0;
wire  [15:0] IN_482_out0;
wire  [15:0] IN_586_out0;
wire  [15:0] IREXEC1_172_out0;
wire  [15:0] IREXEC1_484_out0;
wire  [15:0] IREXEC2_562_out0;
wire  [15:0] IREXEC2_590_out0;
wire  [15:0] IR_22_out0;
wire  [15:0] IR_241_out0;
wire  [15:0] IR_606_out0;
wire  [15:0] MUX1_103_out0;
wire  [15:0] MUX1_192_out0;
wire  [15:0] MUX1_267_out0;
wire  [15:0] MUX1_363_out0;
wire  [15:0] MUX1_408_out0;
wire  [15:0] MUX1_474_out0;
wire  [15:0] MUX1_512_out0;
wire  [15:0] MUX1_54_out0;
wire  [15:0] MUX1_56_out0;
wire  [15:0] MUX1_609_out0;
wire  [15:0] MUX1_630_out0;
wire  [15:0] MUX2_210_out0;
wire  [15:0] MUX2_311_out0;
wire  [15:0] MUX2_324_out0;
wire  [15:0] MUX2_460_out0;
wire  [15:0] MUX3_340_out0;
wire  [15:0] MUX3_40_out0;
wire  [15:0] MUX4_136_out0;
wire  [15:0] MUX4_152_out0;
wire  [15:0] MUX4_231_out0;
wire  [15:0] MUX4_348_out0;
wire  [15:0] MUX4_3_out0;
wire  [15:0] MUX4_469_out0;
wire  [15:0] MUX4_46_out0;
wire  [15:0] MUX4_515_out0;
wire  [15:0] MUX4_576_out0;
wire  [15:0] MUX5_288_out0;
wire  [15:0] MUX5_443_out0;
wire  [15:0] MUX6_169_out0;
wire  [15:0] MUX7_161_out0;
wire  [15:0] MUX7_415_out0;
wire  [15:0] MUX7_589_out0;
wire  [15:0] MUX7_91_out0;
wire  [15:0] N_134_out0;
wire  [15:0] OP1_466_out0;
wire  [15:0] OP1_504_out0;
wire  [15:0] OP2_313_out0;
wire  [15:0] OP2_428_out0;
wire  [15:0] OP2_486_out0;
wire  [15:0] OP2_615_out0;
wire  [15:0] OP2_626_out0;
wire  [15:0] OUT_104_out0;
wire  [15:0] OUT_289_out0;
wire  [15:0] OUT_295_out0;
wire  [15:0] OUT_378_out0;
wire  [15:0] OUT_591_out0;
wire  [15:0] OUT_600_out0;
wire  [15:0] OUT_634_out0;
wire  [15:0] R0TEST_273_out0;
wire  [15:0] R0TEST_370_out0;
wire  [15:0] R0_110_out0;
wire  [15:0] R0_217_out0;
wire  [15:0] R0_595_out0;
wire  [15:0] R1TEST_496_out0;
wire  [15:0] R1TEST_500_out0;
wire  [15:0] R1_416_out0;
wire  [15:0] R1_425_out0;
wire  [15:0] R1_580_out0;
wire  [15:0] R2TEST_524_out0;
wire  [15:0] R2TEST_546_out0;
wire  [15:0] R2_101_out0;
wire  [15:0] R2_256_out0;
wire  [15:0] R2_479_out0;
wire  [15:0] R3TEST_236_out0;
wire  [15:0] R3TEST_24_out0;
wire  [15:0] R3_268_out0;
wire  [15:0] R3_327_out0;
wire  [15:0] R3_433_out0;
wire  [15:0] RAM1_249_out0;
wire  [15:0] RAMDOUT_252_out0;
wire  [15:0] RAMDOUT_5_out0;
wire  [15:0] RDOUT_223_out0;
wire  [15:0] RD_68_out0;
wire  [15:0] REGDIN_551_out0;
wire  [15:0] RM_316_out0;
wire  [15:0] RM_395_out0;
wire  [15:0] RM_541_out0;
wire  [15:0] TESTVIEW_97_out0;
wire  [15:0] XOR1_523_out0;
wire  [15:0] Y_12_out0;
wire  [15:0] Y_599_out0;
wire  [15:0] v_100_out0;
wire  [15:0] v_123_out0;
wire  [15:0] v_186_out0;
wire  [15:0] v_30_out0;
wire  [15:0] v_334_out0;
wire  [15:0] v_342_out0;
wire  [15:0] v_376_out0;
wire  [15:0] v_384_out0;
wire  [15:0] v_388_out0;
wire  [15:0] v_398_out0;
wire  [15:0] v_411_out0;
wire  [15:0] v_423_out0;
wire  [15:0] v_483_out0;
wire  [15:0] v_497_out0;
wire  [15:0] v_528_out0;
wire  [15:0] v_532_out0;
wire  [15:0] v_534_out0;
wire  [15:0] v_572_out0;
wire  [15:0] v_617_out0;
wire  [15:0] v_7_out0;
wire  [1:0] A1_571_out0;
wire  [1:0] AD1_639_out0;
wire  [1:0] AD2_521_out0;
wire  [1:0] AD3_494_out0;
wire  [1:0] C1_527_out0;
wire  [1:0] C1_635_out0;
wire  [1:0] C2_359_out0;
wire  [1:0] C2_475_out0;
wire  [1:0] C3_437_out0;
wire  [1:0] C3_452_out0;
wire  [1:0] D_148_out0;
wire  [1:0] IN0_409_out0;
wire  [1:0] IN15_95_out0;
wire  [1:0] MUX1_167_out0;
wire  [1:0] MUX1_174_out0;
wire  [1:0] MUX2_625_out0;
wire  [1:0] MUX2_90_out0;
wire  [1:0] MUX6_502_out0;
wire  [1:0] M_405_out0;
wire  [1:0] SHIFT_112_out0;
wire  [1:0] SHIFT_213_out0;
wire  [1:0] SHIFT_260_out0;
wire  [1:0] SR_291_out0;
wire  [1:0] SR_32_out0;
wire  [1:0] SR_429_out0;
wire  [1:0] SR_478_out0;
wire  [1:0] v_198_out0;
wire  [1:0] v_25_out1;
wire  [1:0] v_339_out0;
wire  [1:0] v_396_out0;
wire  [1:0] v_414_out0;
wire  [1:0] v_531_out0;
wire  [1:0] v_563_out0;
wire  [2:0] IR1315_245_out0;
wire  [2:0] OP_537_out0;
wire  [2:0] OP_60_out0;
wire  [2:0] OP_84_out0;
wire  [2:0] v_237_out0;
wire  [2:0] v_2_out0;
wire  [2:0] v_317_out0;
wire  [2:0] v_603_out0;
wire  [2:0] v_628_out0;
wire  [3:0] B_355_out0;
wire  [3:0] B_404_out0;
wire  [3:0] C1_88_out0;
wire  [3:0] C2_26_out0;
wire  [3:0] C3_170_out0;
wire  [3:0] IN0_61_out0;
wire  [3:0] IN15_356_out0;
wire  [3:0] MUX2_159_out0;
wire  [3:0] MUX6_154_out0;
wire  [3:0] v_250_out0;
wire  [3:0] v_278_out0;
wire  [3:0] v_300_out0;
wire  [3:0] v_320_out1;
wire  [3:0] v_451_out0;
wire  [3:0] v_489_out0;
wire  [3:0] v_592_out0;
wire  [3:0] v_632_out0;
wire  [4:0] K_16_out0;
wire  [4:0] v_229_out0;
wire  [4:0] v_34_out0;
wire  [4:0] v_417_out0;
wire  [5:0] v_514_out0;
wire  [5:0] v_539_out0;
wire  [6:0] v_397_out0;
wire  [6:0] v_511_out0;
wire  [7:0] C1_263_out0;
wire  [7:0] C1_335_out0;
wire  [7:0] C1_508_out0;
wire  [7:0] C1_593_out0;
wire  [7:0] C1_63_out0;
wire  [7:0] C2_386_out0;
wire  [7:0] IN0_614_out0;
wire  [7:0] IN14_47_out0;
wire  [7:0] IN15_157_out0;
wire  [7:0] IN1_39_out0;
wire  [7:0] MUX1_83_out0;
wire  [7:0] MUX2_243_out0;
wire  [7:0] MUX6_232_out0;
wire  [7:0] v_106_out0;
wire  [7:0] v_162_out0;
wire  [7:0] v_162_out1;
wire  [7:0] v_219_out0;
wire  [7:0] v_281_out0;
wire  [7:0] v_284_out0;
wire  [7:0] v_284_out1;
wire  [7:0] v_347_out0;
wire  [7:0] v_43_out0;
wire  [8:0] C4_298_out0;
wire  [8:0] v_122_out0;
wire  [8:0] v_234_out0;
wire  [9:0] v_332_out0;
wire  [9:0] v_426_out0;
wire A1_225_out1;
wire A1_407_out1;
wire A1_571_out1;
wire A1_597_out1;
wire A1_8_out1;
wire ADC_283_out0;
wire ADC_491_out0;
wire ADD_559_out0;
wire ADD_92_out0;
wire AND_181_out0;
wire AND_296_out0;
wire BIC_353_out0;
wire BIC_570_out0;
wire B_421_out0;
wire B_533_out0;
wire C1_357_out0;
wire C1_390_out0;
wire C1_548_out0;
wire C1_629_out0;
wire C2_228_out0;
wire CALU_380_out0;
wire CALU_509_out0;
wire CALU_552_out0;
wire CFF_11_out0;
wire CMP_393_out0;
wire CMP_6_out0;
wire COUT2_129_out0;
wire COUT_132_out0;
wire COUT_179_out0;
wire COUT_1_out0;
wire COUT_266_out0;
wire COUT_304_out0;
wire COUT_341_out0;
wire COUT_529_out0;
wire COUT_565_out0;
wire C_108_out0;
wire C_109_out0;
wire C_80_out0;
wire D1_445_out0;
wire D1_445_out1;
wire D1_445_out2;
wire D1_445_out3;
wire EN_206_out0;
wire EN_208_out0;
wire EN_211_out0;
wire EN_467_out0;
wire EQ10_73_out0;
wire EQ11_640_out0;
wire EQ1_113_out0;
wire EQ1_137_out0;
wire EQ1_214_out0;
wire EQ1_307_out0;
wire EQ1_389_out0;
wire EQ1_422_out0;
wire EQ1_446_out0;
wire EQ1_535_out0;
wire EQ1_601_out0;
wire EQ2_153_out0;
wire EQ2_185_out0;
wire EQ2_193_out0;
wire EQ2_207_out0;
wire EQ2_258_out0;
wire EQ2_424_out0;
wire EQ3_368_out0;
wire EQ3_471_out0;
wire EQ3_94_out0;
wire EQ4_292_out0;
wire EQ4_35_out0;
wire EQ4_87_out0;
wire EQ5_187_out0;
wire EQ5_277_out0;
wire EQ5_498_out0;
wire EQ6_325_out0;
wire EQ6_382_out0;
wire EQ6_59_out0;
wire EQ7_555_out0;
wire EQ7_624_out0;
wire EQ8_259_out0;
wire EQ9_86_out0;
wire EQ_130_out0;
wire EQ_197_out0;
wire EQ_21_out0;
wire EQ_276_out0;
wire EQ_399_out0;
wire EXEC1_131_out0;
wire EXEC1_149_out0;
wire EXEC1_270_out0;
wire EXEC1_271_out0;
wire EXEC1_530_out0;
wire EXEC1_575_out0;
wire EXEC2_13_out0;
wire EXEC2_209_out0;
wire EXEC2_269_out0;
wire FETCH_119_out0;
wire FETCH_462_out0;
wire G10_31_out0;
wire G10_444_out0;
wire G10_605_out0;
wire G11_17_out0;
wire G11_184_out0;
wire G11_619_out0;
wire G12_216_out0;
wire G12_468_out0;
wire G13_116_out0;
wire G13_15_out0;
wire G14_221_out0;
wire G14_540_out0;
wire G15_351_out0;
wire G15_518_out0;
wire G16_314_out0;
wire G16_98_out0;
wire G1_124_out0;
wire G1_387_out0;
wire G1_413_out0;
wire G1_440_out0;
wire G1_457_out0;
wire G1_513_out0;
wire G1_560_out0;
wire G1_577_out0;
wire G1_622_out0;
wire G1_62_out0;
wire G1_631_out0;
wire G2_175_out0;
wire G2_282_out0;
wire G2_322_out0;
wire G2_542_out0;
wire G2_549_out0;
wire G2_567_out0;
wire G2_620_out0;
wire G2_627_out0;
wire G2_81_out0;
wire G3_133_out0;
wire G3_235_out0;
wire G3_29_out0;
wire G3_379_out0;
wire G3_506_out0;
wire G3_582_out0;
wire G4_147_out0;
wire G4_321_out0;
wire G4_371_out0;
wire G4_373_out0;
wire G4_558_out0;
wire G5_195_out0;
wire G5_253_out0;
wire G5_344_out0;
wire G5_402_out0;
wire G5_472_out0;
wire G6_120_out0;
wire G6_255_out0;
wire G6_346_out0;
wire G6_545_out0;
wire G6_556_out0;
wire G6_66_out0;
wire G7_218_out0;
wire G7_230_out0;
wire G7_449_out0;
wire G7_536_out0;
wire G7_573_out0;
wire G8_328_out0;
wire G8_337_out0;
wire G8_430_out0;
wire G8_463_out0;
wire G8_470_out0;
wire G8_583_out0;
wire G9_191_out0;
wire G9_212_out0;
wire G9_406_out0;
wire G9_578_out0;
wire G9_57_out0;
wire IN0_28_out0;
wire IN15_121_out0;
wire IR15_183_out0;
wire IR15_326_out0;
wire JEQN_4_out0;
wire JEQ_643_out0;
wire JMIN_64_out0;
wire JMI_0_out0;
wire JMPN_242_out0;
wire JMP_82_out0;
wire LDSTB_434_out0;
wire LDSTB_53_out0;
wire LDST_301_out0;
wire LDST_381_out0;
wire L_427_out0;
wire MI_142_out0;
wire MI_201_out0;
wire MI_37_out0;
wire MI_76_out0;
wire MI_93_out0;
wire MOV_168_out0;
wire MOV_394_out0;
wire MUX2_280_out0;
wire MUX2_455_out0;
wire MUX3_436_out0;
wire MUX6_9_out0;
wire MVN_248_out0;
wire MVN_448_out0;
wire P_67_out0;
wire RAMWEN_44_out0;
wire RAMWEN_522_out0;
wire SBC_202_out0;
wire SBC_23_out0;
wire STALL0_177_out0;
wire STALL0_188_out0;
wire STALL0_233_out0;
wire STALL0_525_out0;
wire STALL0_612_out0;
wire STALLE1_308_out0;
wire STALLE1_345_out0;
wire STALLE1_365_out0;
wire STALLE1_375_out0;
wire STALLE1_505_out0;
wire STALLE2_140_out0;
wire STALLE2_144_out0;
wire STALLE2_55_out0;
wire STALLF_244_out0;
wire STALLF_310_out0;
wire STALLF_516_out0;
wire STALLF_70_out0;
wire STALLF_71_out0;
wire STALLF_77_out0;
wire STP_400_out0;
wire STP_473_out0;
wire SUB_146_out0;
wire SUB_438_out0;
wire S_14_out0;
wire S_377_out0;
wire S_453_out0;
wire TST_336_out0;
wire TST_611_out0;
wire U_126_out0;
wire WENALU_141_out0;
wire WENALU_303_out0;
wire WENALU_585_out0;
wire WENALU_636_out0;
wire WENLDST_633_out0;
wire WENRAM_166_out0;
wire WREN3_111_out0;
wire W_254_out0;
wire v_105_out0;
wire v_114_out0;
wire v_117_out0;
wire v_125_out0;
wire v_135_out0;
wire v_155_out0;
wire v_158_out0;
wire v_165_out0;
wire v_178_out0;
wire v_180_out0;
wire v_194_out0;
wire v_196_out0;
wire v_199_out0;
wire v_19_out0;
wire v_215_out0;
wire v_220_out0;
wire v_224_out0;
wire v_226_out0;
wire v_226_out1;
wire v_227_out0;
wire v_238_out0;
wire v_239_out0;
wire v_247_out0;
wire v_264_out0;
wire v_27_out0;
wire v_286_out0;
wire v_287_out0;
wire v_290_out0;
wire v_293_out0;
wire v_294_out0;
wire v_299_out0;
wire v_302_out0;
wire v_309_out0;
wire v_312_out0;
wire v_318_out0;
wire v_323_out0;
wire v_329_out0;
wire v_331_out0;
wire v_338_out0;
wire v_33_out0;
wire v_354_out0;
wire v_360_out0;
wire v_362_out0;
wire v_364_out0;
wire v_364_out1;
wire v_36_out0;
wire v_374_out0;
wire v_383_out0;
wire v_385_out0;
wire v_391_out0;
wire v_435_out0;
wire v_439_out0;
wire v_441_out0;
wire v_447_out0;
wire v_45_out0;
wire v_480_out0;
wire v_481_out0;
wire v_485_out0;
wire v_487_out0;
wire v_492_out0;
wire v_495_out0;
wire v_501_out0;
wire v_507_out0;
wire v_517_out0;
wire v_519_out0;
wire v_526_out0;
wire v_52_out1;
wire v_561_out0;
wire v_574_out0;
wire v_581_out0;
wire v_594_out0;
wire v_596_out0;
wire v_598_out0;
wire v_602_out0;
wire v_604_out0;
wire v_616_out0;
wire v_638_out0;
wire v_72_out0;
wire v_75_out0;
wire v_78_out0;
wire v_85_out0;
wire v_96_out0;
wire v_99_out0;

always @(posedge clk) REG1_50_out0 <= EXEC1_270_out0 ? DIN_203_out0 : REG1_50_out0;
always @(posedge clk) REG1_51_out0 <= EXEC1_271_out0 ? DIN_204_out0 : REG1_51_out0;
always @(posedge clk) FF2_128_out0 <= FF1_459_out0;
always @(posedge clk) REG1_156_out0 <= G1_124_out0 ? A1_571_out0 : REG1_156_out0;
always @(posedge clk) REG1_164_out0 <= D1_445_out1 ? DIN3_461_out0 : REG1_164_out0;
RAM1_249 I1 (RAM1_249_out0, MUX1_392_out0, RDOUT_223_out0, RAMWEN_44_out0, clk);
always @(posedge clk) FF1_251_out0 <= G5_344_out0 ? G4_373_out0 : FF1_251_out0;
always @(posedge clk) REG1_274_out0 <= MUX2_455_out0 ? MUX1_272_out0 : REG1_274_out0;
always @(posedge clk) REG3_333_out0 <= D1_445_out3 ? DIN3_461_out0 : REG3_333_out0;
always @(posedge clk) Z_361_out0 <= EXEC2_209_out0 ? COUT_304_out0 : Z_361_out0;
always @(posedge clk) FF1_459_out0 <= G2_620_out0;
always @(posedge clk) FF1_538_out0 <= G2_567_out0 ? CFF_11_out0 : FF1_538_out0;
always @(posedge clk) REG0_543_out0 <= D1_445_out0 ? DIN3_461_out0 : REG0_543_out0;
always @(posedge clk) N_564_out0 <= EXEC2_209_out0 ? EQ1_446_out0 : N_564_out0;
always @(posedge clk) REG2_584_out0 <= D1_445_out2 ? DIN3_461_out0 : REG2_584_out0;
always @(posedge clk) FF2_621_out0 <= C1_629_out0;
assign C1_635_out0 = 2'h0;
assign C1_629_out0 = 1'h1;
assign C1_593_out0 = 8'h0;
assign C2_579_out0 = 12'hfff;
assign C2_550_out0 = 12'h1;
assign C1_548_out0 = 1'h0;
assign C1_544_out0 = 16'hffff;
assign C1_527_out0 = 2'h3;
assign C1_508_out0 = 8'h0;
assign C2_475_out0 = 2'h1;
assign C3_452_out0 = 2'h0;
assign C3_437_out0 = 2'h2;
assign C3_431_out0 = 12'h1;
assign C1_390_out0 = 1'h0;
assign C2_386_out0 = 8'hff;
assign C1_367_out0 = 11'h0;
assign C2_359_out0 = 2'h3;
assign C1_357_out0 = 1'h0;
assign C1_335_out0 = 8'h0;
assign C4_298_out0 = 9'h0;
assign C1_263_out0 = 8'h0;
assign C2_228_out0 = 1'h0;
assign C3_170_out0 = 4'h0;
assign C1_88_out0 = 4'h0;
assign C1_63_out0 = 8'h0;
assign C2_26_out0 = 4'hff;
assign COUT_1_out0 = FF1_538_out0;
assign EXEC2_13_out0 = FF2_128_out0;
assign EQ_21_out0 = Z_361_out0;
assign C_80_out0 = FF1_538_out0;
assign R0_110_out0 = REG0_543_out0;
assign DOUT_138_out0 = REG1_50_out0;
assign DOUT_139_out0 = REG1_51_out0;
assign DIN_173_out0 = RAM1_249_out0;
assign MI_201_out0 = N_564_out0;
assign EQ2_207_out0 = REG1_156_out0 == 2'h2;
assign {A1_225_out1,A1_225_out0 } = REG1_274_out0 + C2_550_out0 + C1_548_out0;
assign RAMDOUT_252_out0 = RAM1_249_out0;
assign R2_256_out0 = REG2_584_out0;
assign RAMOUT_262_out0 = RAM1_249_out0;
assign R3_327_out0 = REG3_333_out0;
assign EQ3_368_out0 = REG1_156_out0 == 2'h0;
assign G4_373_out0 = ! FF1_251_out0;
assign EQ1_422_out0 = REG1_156_out0 == 2'h1;
assign R1_425_out0 = REG1_164_out0;
assign EXEC1_575_out0 = FF1_459_out0;
assign PCOUT_637_out0 = REG1_274_out0;
assign RAMDOUT_5_out0 = RAMDOUT_252_out0;
assign STALLE2_55_out0 = EQ2_207_out0;
assign MI_76_out0 = MI_201_out0;
assign COUT_132_out0 = A1_225_out1;
assign EXEC1_149_out0 = EXEC1_575_out0;
assign IREXEC1_172_out0 = DOUT_138_out0;
assign MUX1_174_out0 = EQ2_207_out0 ? C3_437_out0 : C2_475_out0;
assign COUT_179_out0 = COUT_1_out0;
assign EQ_197_out0 = EQ_21_out0;
assign R3TEST_236_out0 = R3_327_out0;
assign MUX1_267_out0 = G4_373_out0 ? DOUT_139_out0 : DOUT_138_out0;
assign EXEC2_269_out0 = EXEC2_13_out0;
assign R0TEST_273_out0 = R0_110_out0;
assign COUT_304_out0 = COUT_1_out0;
assign STALLE1_308_out0 = EQ1_422_out0;
assign R1TEST_496_out0 = R1_425_out0;
assign DM1_510_out0 = FF1_251_out0 ? 16'h0 : DIN_173_out0;
assign DM1_510_out1 = FF1_251_out0 ? DIN_173_out0 : 16'h0;
assign R2TEST_524_out0 = R2_256_out0;
assign CALU_552_out0 = COUT_1_out0;
assign IREXEC2_590_out0 = DOUT_139_out0;
assign STALL0_612_out0 = EQ3_368_out0;
assign R3TEST_24_out0 = R3TEST_236_out0;
assign MI_37_out0 = MI_76_out0;
assign EXEC1_131_out0 = EXEC1_149_out0;
assign STALLE2_144_out0 = STALLE2_55_out0;
assign STALL0_177_out0 = STALL0_612_out0;
assign DIN_203_out0 = DM1_510_out0;
assign DIN_204_out0 = DM1_510_out1;
assign EXEC2_209_out0 = EXEC2_269_out0;
assign MUX2_210_out0 = FF2_621_out0 ? MUX1_267_out0 : DIN_173_out0;
assign EQ_276_out0 = EQ_197_out0;
assign v_347_out0 = RAMDOUT_5_out0[7:0];
assign STALLE1_365_out0 = STALLE1_308_out0;
assign R0TEST_370_out0 = R0TEST_273_out0;
assign IREXEC1_484_out0 = IREXEC1_172_out0;
assign R1TEST_500_out0 = R1TEST_496_out0;
assign CALU_509_out0 = CALU_552_out0;
assign COUT_529_out0 = COUT_179_out0;
assign EXEC1_530_out0 = EXEC1_149_out0;
assign R2TEST_546_out0 = R2TEST_524_out0;
assign IREXEC2_562_out0 = IREXEC2_590_out0;
assign {A1_571_out1,A1_571_out0 } = REG1_156_out0 + MUX1_174_out0 + C1_390_out0;
assign G3_29_out0 = ! STALLE1_365_out0;
assign MI_93_out0 = MI_37_out0;
assign R2_101_out0 = R2TEST_546_out0;
assign v_123_out0 = { v_347_out0,C1_335_out0 };
assign EQ_130_out0 = EQ_276_out0;
assign N_134_out0 = MUX2_210_out0;
assign STALLE2_140_out0 = STALLE2_144_out0;
assign MI_142_out0 = MI_37_out0;
assign R0_217_out0 = R0TEST_370_out0;
assign STALLE1_345_out0 = STALLE1_365_out0;
assign IROUT_350_out0 = IREXEC1_484_out0;
assign CALU_380_out0 = CALU_509_out0;
assign EQ_399_out0 = EQ_276_out0;
assign R3_433_out0 = R3TEST_24_out0;
assign STALL0_525_out0 = STALL0_177_out0;
assign COUT_565_out0 = A1_571_out1;
assign R1_580_out0 = R1TEST_500_out0;
assign v_592_out0 = MUX2_210_out0[15:12];
assign EQ6_59_out0 = v_592_out0 == 4'h2;
assign EQ10_73_out0 = v_592_out0 == 4'h9;
assign EQ9_86_out0 = v_592_out0 == 4'h8;
assign EQ4_87_out0 = v_592_out0 == 4'hb;
assign EQ3_94_out0 = v_592_out0 == 4'hd;
assign v_102_out0 = N_134_out0[11:0];
assign EQ2_185_out0 = v_592_out0 == 4'hc;
assign EQ5_187_out0 = v_592_out0 == 4'h4;
assign STALL0_188_out0 = STALL0_525_out0;
assign G9_191_out0 = G4_373_out0 && G3_29_out0;
assign EQ1_214_out0 = v_592_out0 == 4'h1;
assign G7_230_out0 = FF1_251_out0 && G3_29_out0;
assign IR_241_out0 = N_134_out0;
assign EQ8_259_out0 = v_592_out0 == 4'h7;
assign R3_268_out0 = R3_433_out0;
assign EQ4_292_out0 = v_592_out0 == 4'he;
assign EQ1_307_out0 = v_592_out0 == 4'h0;
assign EQ6_325_out0 = v_592_out0 == 4'h5;
assign STALLE1_375_out0 = STALLE1_345_out0;
assign R1_416_out0 = R1_580_out0;
assign R2_479_out0 = R2_101_out0;
assign EQ5_498_out0 = v_592_out0 == 4'hf;
assign EQ7_555_out0 = v_592_out0 == 4'h6;
assign R0_595_out0 = R0_217_out0;
assign EQ7_624_out0 = v_592_out0 == 4'h3;
assign EQ11_640_out0 = v_592_out0 == 4'ha;
assign v_2_out0 = IR_241_out0[14:12];
assign JEQN_4_out0 = EQ7_555_out0;
assign SBC_23_out0 = EQ4_87_out0;
assign R0OUT_38_out0 = R0_595_out0;
assign R1OUT_49_out0 = R1_416_out0;
assign LDSTB_53_out0 = EQ1_214_out0;
assign JMIN_64_out0 = EQ6_325_out0;
assign G6_120_out0 = MI_93_out0 && EQ6_325_out0;
assign R3OUT_127_out0 = R3_268_out0;
assign SUB_146_out0 = EQ10_73_out0;
assign R2OUT_163_out0 = R2_479_out0;
assign G2_175_out0 = EQ_130_out0 && EQ7_555_out0;
assign v_198_out0 = IR_241_out0[1:0];
assign STALL0_233_out0 = STALL0_188_out0;
assign JMPN_242_out0 = EQ5_187_out0;
assign EXEC1_270_out0 = G9_191_out0;
assign EXEC1_271_out0 = G7_230_out0;
assign AND_296_out0 = EQ4_292_out0;
assign LDST_301_out0 = EQ1_307_out0;
assign TST_336_out0 = EQ5_498_out0;
assign STALL0_352_out0 = STALL0_188_out0;
assign v_385_out0 = IR_241_out0[15:15];
assign CMP_393_out0 = EQ3_94_out0;
assign MOV_394_out0 = EQ2_185_out0;
assign STP_400_out0 = EQ8_259_out0;
assign G10_444_out0 = EQ1_307_out0 || EQ1_214_out0;
assign MVN_448_out0 = EQ7_624_out0;
assign ADC_491_out0 = EQ11_640_out0;
assign STALLE1_505_out0 = STALLE1_375_out0;
assign v_531_out0 = IR_241_out0[11:10];
assign ADD_559_out0 = EQ9_86_out0;
assign v_561_out0 = IR_241_out0[5:5];
assign BIC_570_out0 = EQ6_59_out0;
assign N_587_out0 = v_102_out0;
assign v_602_out0 = IR_241_out0[12:12];
assign IR_606_out0 = IR_241_out0;
assign JMI_0_out0 = JMIN_64_out0;
assign CMP_6_out0 = CMP_393_out0;
assign S_14_out0 = v_561_out0;
assign IR_22_out0 = IR_606_out0;
assign JMP_82_out0 = JMPN_242_out0;
assign OP_84_out0 = v_2_out0;
assign ADD_92_out0 = ADD_559_out0;
assign D_148_out0 = v_531_out0;
assign MOV_168_out0 = MOV_394_out0;
assign v_178_out0 = IR_606_out0[8:8];
assign AND_181_out0 = AND_296_out0;
assign IR15_183_out0 = v_385_out0;
assign SBC_202_out0 = SBC_23_out0;
assign v_229_out0 = IR_606_out0[4:0];
assign MVN_248_out0 = MVN_448_out0;
assign ADC_283_out0 = ADC_491_out0;
assign v_300_out0 = IR_606_out0[7:4];
assign v_338_out0 = IR_606_out0[9:9];
assign BIC_353_out0 = BIC_570_out0;
assign LDST_381_out0 = LDST_301_out0;
assign M_405_out0 = v_198_out0;
assign B_421_out0 = v_602_out0;
assign LDSTB_434_out0 = LDSTB_53_out0;
assign SUB_438_out0 = SUB_146_out0;
assign STP_473_out0 = STP_400_out0;
assign v_563_out0 = IR_606_out0[3:2];
assign G8_583_out0 = G2_175_out0 || G6_120_out0;
assign TST_611_out0 = TST_336_out0;
assign JEQ_643_out0 = JEQN_4_out0;
assign K_16_out0 = v_229_out0;
assign OP_60_out0 = OP_84_out0;
assign v_85_out0 = IR_22_out0[5:5];
assign MUX2_90_out0 = EXEC2_269_out0 ? D_148_out0 : M_405_out0;
assign C_108_out0 = v_338_out0;
assign EQ1_113_out0 = OP_84_out0 == 3'h2;
assign EQ2_153_out0 = OP_84_out0 == 3'h3;
assign v_155_out0 = IR_22_out0[7:7];
assign v_237_out0 = IR_22_out0[4:2];
assign v_247_out0 = IR_22_out0[6:6];
assign G6_255_out0 = MI_142_out0 && JMI_0_out0;
assign SHIFT_260_out0 = v_563_out0;
assign IR15_326_out0 = IR15_183_out0;
assign S_377_out0 = v_178_out0;
assign v_391_out0 = IR_22_out0[12:12];
assign B_404_out0 = v_300_out0;
assign G1_413_out0 = EQ_399_out0 && JEQ_643_out0;
assign v_451_out0 = IR_22_out0[5:2];
assign v_481_out0 = IR_22_out0[8:8];
assign G1_513_out0 = G10_444_out0 || G8_583_out0;
assign AD2_521_out0 = M_405_out0;
assign G2_549_out0 = ! STP_473_out0;
assign v_594_out0 = IR_22_out0[9:9];
assign v_628_out0 = IR_22_out0[15:13];
assign AD1_639_out0 = D_148_out0;
assign G11_17_out0 = FF2_621_out0 && G1_513_out0;
assign EQ4_35_out0 = OP_60_out0 == 3'h5;
assign P_67_out0 = v_155_out0;
assign v_89_out0 = { v_451_out0,C1_508_out0 };
assign C_109_out0 = C_108_out0;
assign SHIFT_112_out0 = SHIFT_260_out0;
assign U_126_out0 = v_247_out0;
assign v_226_out0 = AD2_521_out0[0:0];
assign v_226_out1 = AD2_521_out0[1:1];
assign IR1315_245_out0 = v_628_out0;
assign W_254_out0 = v_481_out0;
assign EQ2_258_out0 = OP_60_out0 == 3'h6;
assign EQ5_277_out0 = OP_60_out0 == 3'h2;
assign B_355_out0 = B_404_out0;
assign v_364_out0 = AD1_639_out0[0:0];
assign v_364_out1 = AD1_639_out0[1:1];
assign EQ6_382_out0 = OP_60_out0 == 3'h3;
assign L_427_out0 = v_594_out0;
assign G8_430_out0 = G1_413_out0 || G6_255_out0;
assign S_453_out0 = v_85_out0;
assign G1_457_out0 = EQ1_113_out0 || EQ2_153_out0;
assign EQ3_471_out0 = OP_60_out0 == 3'h7;
assign AD3_494_out0 = MUX2_90_out0;
assign v_499_out0 = { v_237_out0,C4_298_out0 };
assign v_528_out0 = { K_16_out0,C1_367_out0 };
assign B_533_out0 = v_391_out0;
assign EQ1_535_out0 = OP_60_out0 == 3'h4;
assign OP_537_out0 = OP_60_out0;
assign G2_567_out0 = S_377_out0 && EXEC1_530_out0;
assign v_36_out0 = B_355_out0[2:2];
assign MUX4_46_out0 = v_226_out0 ? R1_425_out0 : R0_110_out0;
assign G9_57_out0 = G8_430_out0 || JMP_82_out0;
assign G6_66_out0 = EQ5_277_out0 || EQ6_382_out0;
assign v_72_out0 = OP_537_out0[1:1];
assign G3_133_out0 = EQ2_258_out0 || EQ3_471_out0;
assign MUX1_167_out0 = C_109_out0 ? C1_527_out0 : SHIFT_112_out0;
assign MUX1_192_out0 = v_364_out0 ? REG1_164_out0 : REG0_543_out0;
assign EQ2_193_out0 = IR1315_245_out0 == 3'h0;
assign G5_195_out0 = B_533_out0 && S_453_out0;
assign SHIFT_213_out0 = SHIFT_112_out0;
assign G7_218_out0 = ! L_427_out0;
assign v_220_out0 = OP_537_out0[0:0];
assign v_238_out0 = B_355_out0[0:0];
assign STALLF_310_out0 = G11_17_out0;
assign MUX2_324_out0 = v_364_out0 ? REG3_333_out0 : REG2_584_out0;
assign MUX4_348_out0 = B_533_out0 ? v_123_out0 : RAMDOUT_5_out0;
assign v_374_out0 = B_355_out0[1:1];
assign G3_379_out0 = ! U_126_out0;
assign EQ1_389_out0 = B_355_out0 == 4'h0;
assign MUX5_443_out0 = v_226_out0 ? R3_327_out0 : R2_256_out0;
assign MUX5_458_out0 = B_533_out0 ? v_499_out0 : v_89_out0;
assign G2_542_out0 = IR15_183_out0 || G1_457_out0;
assign G6_545_out0 = W_254_out0 && EXEC1_131_out0;
assign G4_558_out0 = !(EQ3_471_out0 || EQ4_35_out0);
assign G1_577_out0 = ! C_109_out0;
assign v_604_out0 = B_355_out0[3:3];
assign SR_32_out0 = MUX1_167_out0;
assign MUX3_40_out0 = v_364_out1 ? MUX2_324_out0 : MUX1_192_out0;
assign STALLF_70_out0 = STALLF_310_out0;
assign G2_81_out0 = G1_577_out0 && v_238_out0;
assign EQ1_137_out0 = SHIFT_213_out0 == 2'h0;
assign MUX6_169_out0 = v_226_out1 ? MUX5_443_out0 : MUX4_46_out0;
assign EN_206_out0 = v_604_out0;
assign EN_208_out0 = v_374_out0;
assign G3_235_out0 = G1_577_out0 && EQ1_389_out0;
assign MUX1_272_out0 = G9_57_out0 ? N_587_out0 : A1_225_out0;
assign MUX2_280_out0 = v_72_out0 ? C_80_out0 : v_220_out0;
assign SR_291_out0 = MUX1_167_out0;
assign G5_344_out0 = !(STALLF_310_out0 && STALL0_177_out0);
assign G1_387_out0 = G6_545_out0 || EXEC2_209_out0;
assign EQ2_424_out0 = SHIFT_213_out0 == 2'h2;
assign SR_429_out0 = MUX1_167_out0;
assign N_456_out0 = MUX5_458_out0;
assign EN_467_out0 = v_36_out0;
assign G8_470_out0 = G3_133_out0 || G6_66_out0;
assign SR_478_out0 = MUX1_167_out0;
assign STALLF_516_out0 = STALLF_310_out0;
assign G7_573_out0 = G6_66_out0 || IR15_326_out0;
assign EQ1_601_out0 = SHIFT_213_out0 == 2'h3;
assign G2_627_out0 = G7_218_out0 && EXEC2_209_out0;
assign G1_62_out0 = EXEC1_530_out0 && G7_573_out0;
assign STALLF_77_out0 = STALLF_516_out0;
assign v_96_out0 = SR_429_out0[1:1];
assign v_105_out0 = SR_32_out0[1:1];
assign DOUT1_107_out0 = MUX3_40_out0;
assign DOUT2_118_out0 = MUX6_169_out0;
assign G1_124_out0 = STALLF_70_out0 || EQ2_207_out0;
assign G4_147_out0 = G1_387_out0 && L_427_out0;
assign v_158_out0 = SR_478_out0[1:1];
assign v_194_out0 = SR_429_out0[0:0];
assign EN_211_out0 = G2_81_out0;
assign v_290_out0 = SR_478_out0[0:0];
assign v_309_out0 = SR_291_out0[0:0];
assign G8_337_out0 = G2_627_out0 && EQ2_193_out0;
assign v_362_out0 = SR_32_out0[0:0];
assign XOR1_588_out0 = N_456_out0 ^ C2_579_out0;
assign v_598_out0 = SR_291_out0[1:1];
assign G1_631_out0 = EQ1_137_out0 || EQ1_601_out0;
assign v_43_out0 = DOUT1_107_out0[7:0];
assign RD_68_out0 = DOUT1_107_out0;
assign STALLF_71_out0 = STALLF_77_out0;
assign v_106_out0 = DOUT1_107_out0[15:8];
assign STALLF_182_out0 = STALLF_77_out0;
assign MUX3_205_out0 = G3_379_out0 ? XOR1_588_out0 : N_456_out0;
assign STALLF_244_out0 = STALLF_77_out0;
assign RM_395_out0 = DOUT2_118_out0;
assign G5_402_out0 = G1_62_out0 && G4_558_out0;
assign G9_406_out0 = G4_147_out0 && EQ2_193_out0;
assign G1_440_out0 = STALL0_188_out0 && STALLF_77_out0;
assign RAMWEN_522_out0 = G8_337_out0;
assign RM_541_out0 = DOUT2_118_out0;
assign MUX1_83_out0 = S_14_out0 ? v_106_out0 : v_43_out0;
assign WENRAM_166_out0 = RAMWEN_522_out0;
assign RM_316_out0 = RM_395_out0;
assign MUX1_408_out0 = C_108_out0 ? v_528_out0 : RM_541_out0;
assign MUX2_455_out0 = STALLF_244_out0 ? STALLE1_505_out0 : G2_549_out0;
assign OP1_504_out0 = RD_68_out0;
assign G2_620_out0 = !(STALL0_233_out0 && STALLF_71_out0);
assign WENLDST_633_out0 = G9_406_out0;
assign WENALU_636_out0 = G5_402_out0;
assign RAMWEN_44_out0 = WENRAM_166_out0;
assign A_65_out0 = MUX1_408_out0;
assign v_74_out0 = RM_316_out0[11:0];
assign WENALU_141_out0 = WENALU_636_out0;
assign v_250_out0 = RM_316_out0[15:12];
assign v_411_out0 = { MUX1_83_out0,C1_593_out0 };
assign FETCH_462_out0 = G2_620_out0;
assign OP1_466_out0 = OP1_504_out0;
assign A_493_out0 = OP1_504_out0;
assign WENALU_585_out0 = WENALU_636_out0;
assign {A1_8_out1,A1_8_out0 } = v_74_out0 + MUX3_205_out0 + G3_379_out0;
assign v_27_out0 = A_493_out0[13:13];
assign v_33_out0 = A_493_out0[2:2];
assign v_78_out0 = A_493_out0[5:5];
assign v_114_out0 = A_493_out0[11:11];
assign FETCH_119_out0 = FETCH_462_out0;
assign v_135_out0 = A_493_out0[8:8];
assign v_196_out0 = A_493_out0[4:4];
assign v_227_out0 = A_493_out0[3:3];
assign v_239_out0 = A_493_out0[7:7];
assign v_286_out0 = A_493_out0[10:10];
assign v_287_out0 = A_493_out0[15:15];
assign MUX5_288_out0 = B_421_out0 ? v_411_out0 : DOUT1_107_out0;
assign v_302_out0 = A_493_out0[0:0];
assign WENALU_303_out0 = WENALU_585_out0;
assign v_312_out0 = A_493_out0[6:6];
assign IN_358_out0 = A_65_out0;
assign MUX3_436_out0 = G2_542_out0 ? WENALU_141_out0 : WENLDST_633_out0;
assign v_441_out0 = A_493_out0[14:14];
assign v_480_out0 = A_493_out0[1:1];
assign v_517_out0 = A_493_out0[9:9];
assign A_568_out0 = A_65_out0;
assign FETCH_569_out0 = FETCH_462_out0;
assign v_574_out0 = A_493_out0[12:12];
assign v_18_out0 = A_568_out0[15:1];
assign v_42_out0 = A_568_out0[14:0];
assign v_52_out0 = IN_358_out0[14:0];
assign v_52_out1 = IN_358_out0[15:1];
assign WREN3_111_out0 = MUX3_436_out0;
assign RDOUT_223_out0 = MUX5_288_out0;
assign COUT_266_out0 = A1_8_out1;
assign v_293_out0 = IN_358_out0[0:0];
assign v_293_out1 = IN_358_out0[15:15];
assign v_532_out0 = { A1_8_out0,v_250_out0 };
assign MUX2_642_out0 = P_67_out0 ? A1_8_out0 : v_74_out0;
assign IN0_28_out0 = v_293_out0;
assign IN1_41_out0 = v_18_out0;
assign IN15_121_out0 = v_52_out1;
assign MUX1_363_out0 = G6_545_out0 ? v_532_out0 : MUX4_348_out0;
assign {A1_407_out1,A1_407_out0 } = MUX2_642_out0 + C3_431_out0 + C2_228_out0;
assign IN14_442_out0 = v_52_out0;
assign D1_445_out0 = (AD3_494_out0 == 2'b00) ? WREN3_111_out0 : 1'h0;
assign D1_445_out1 = (AD3_494_out0 == 2'b01) ? WREN3_111_out0 : 1'h0;
assign D1_445_out2 = (AD3_494_out0 == 2'b10) ? WREN3_111_out0 : 1'h0;
assign D1_445_out3 = (AD3_494_out0 == 2'b11) ? WREN3_111_out0 : 1'h0;
assign IN1_477_out0 = v_293_out1;
assign IN14_610_out0 = v_42_out0;
assign MUX6_9_out0 = v_309_out0 ? IN0_28_out0 : IN15_121_out0;
assign MUX6_69_out0 = G5_195_out0 ? A1_407_out0 : MUX2_642_out0;
assign COUT2_129_out0 = A1_407_out1;
assign v_398_out0 = { IN1_41_out0,CALU_380_out0 };
assign v_497_out0 = { C1_357_out0,IN14_442_out0 };
assign REGDIN_551_out0 = MUX1_363_out0;
assign v_572_out0 = { IN1_477_out0,C1_357_out0 };
assign v_617_out0 = { CALU_380_out0,IN14_610_out0 };
assign v_7_out0 = { IN1_477_out0,MUX6_9_out0 };
assign MUX4_152_out0 = v_309_out0 ? v_572_out0 : v_497_out0;
assign RAMADDRMUX_160_out0 = MUX6_69_out0;
assign MUX4_576_out0 = EQ2_424_out0 ? v_398_out0 : v_617_out0;
assign RAMADDRMUX_20_out0 = RAMADDRMUX_160_out0;
assign MUX1_103_out0 = G1_631_out0 ? A_568_out0 : MUX4_576_out0;
assign MUX7_161_out0 = v_598_out0 ? v_7_out0 : MUX4_152_out0;
assign MUX1_56_out0 = EN_211_out0 ? MUX7_161_out0 : IN_358_out0;
assign OUT_104_out0 = MUX1_103_out0;
assign MUX1_392_out0 = G1_440_out0 ? RAMADDRMUX_20_out0 : PCOUT_637_out0;
assign OUT_634_out0 = MUX1_56_out0;
assign IN_586_out0 = OUT_634_out0;
assign v_25_out0 = IN_586_out0[13:0];
assign v_25_out1 = IN_586_out0[15:2];
assign v_339_out0 = IN_586_out0[1:0];
assign v_339_out1 = IN_586_out0[15:14];
assign v_439_out0 = IN_586_out0[15:15];
assign IN15_95_out0 = v_25_out1;
assign IN14_189_out0 = v_25_out0;
assign IN1_257_out0 = v_339_out1;
assign IN0_409_out0 = v_339_out0;
assign MUX2_625_out0 = v_439_out0 ? C2_359_out0 : C3_452_out0;
assign v_376_out0 = { C1_635_out0,IN14_189_out0 };
assign v_384_out0 = { IN1_257_out0,C1_635_out0 };
assign MUX6_502_out0 = v_290_out0 ? IN0_409_out0 : MUX2_625_out0;
assign v_186_out0 = { IN1_257_out0,MUX6_502_out0 };
assign MUX4_469_out0 = v_290_out0 ? v_384_out0 : v_376_out0;
assign MUX7_415_out0 = v_158_out0 ? v_186_out0 : MUX4_469_out0;
assign MUX1_630_out0 = EN_208_out0 ? MUX7_415_out0 : IN_586_out0;
assign OUT_289_out0 = MUX1_630_out0;
assign IN_482_out0 = OUT_289_out0;
assign v_320_out0 = IN_482_out0[11:0];
assign v_320_out1 = IN_482_out0[15:4];
assign v_354_out0 = IN_482_out0[15:15];
assign v_489_out0 = IN_482_out0[3:0];
assign v_489_out1 = IN_482_out0[15:12];
assign IN0_61_out0 = v_489_out0;
assign MUX2_159_out0 = v_354_out0 ? C2_26_out0 : C3_170_out0;
assign IN15_356_out0 = v_320_out1;
assign IN14_450_out0 = v_320_out0;
assign IN1_465_out0 = v_489_out1;
assign MUX6_154_out0 = v_194_out0 ? IN0_61_out0 : MUX2_159_out0;
assign v_342_out0 = { IN1_465_out0,C1_88_out0 };
assign v_483_out0 = { C1_88_out0,IN14_450_out0 };
assign v_388_out0 = { IN1_465_out0,MUX6_154_out0 };
assign MUX4_515_out0 = v_194_out0 ? v_342_out0 : v_483_out0;
assign MUX7_91_out0 = v_96_out0 ? v_388_out0 : MUX4_515_out0;
assign MUX1_54_out0 = EN_467_out0 ? MUX7_91_out0 : IN_482_out0;
assign OUT_591_out0 = MUX1_54_out0;
assign IN_143_out0 = OUT_591_out0;
assign v_117_out0 = IN_143_out0[15:15];
assign v_162_out0 = IN_143_out0[7:0];
assign v_162_out1 = IN_143_out0[15:8];
assign v_284_out0 = IN_143_out0[7:0];
assign v_284_out1 = IN_143_out0[15:8];
assign IN1_39_out0 = v_284_out1;
assign IN14_47_out0 = v_162_out0;
assign IN15_157_out0 = v_162_out1;
assign MUX2_243_out0 = v_117_out0 ? C2_386_out0 : C1_263_out0;
assign IN0_614_out0 = v_284_out0;
assign v_30_out0 = { IN1_39_out0,C1_63_out0 };
assign MUX6_232_out0 = v_362_out0 ? IN0_614_out0 : MUX2_243_out0;
assign v_534_out0 = { C1_63_out0,IN14_47_out0 };
assign v_100_out0 = { IN1_39_out0,MUX6_232_out0 };
assign MUX4_136_out0 = v_362_out0 ? v_30_out0 : v_534_out0;
assign MUX7_589_out0 = v_105_out0 ? v_100_out0 : MUX4_136_out0;
assign MUX1_474_out0 = EN_206_out0 ? MUX7_589_out0 : IN_143_out0;
assign OUT_378_out0 = MUX1_474_out0;
assign MUX2_311_out0 = G3_235_out0 ? OUT_104_out0 : OUT_378_out0;
assign OUT_600_out0 = MUX2_311_out0;
assign OP2_313_out0 = OUT_600_out0;
assign OP2_486_out0 = OP2_313_out0;
assign OP2_626_out0 = OP2_313_out0;
assign A_366_out0 = OP2_486_out0;
assign OP2_428_out0 = OP2_626_out0;
assign OP2_615_out0 = OP2_486_out0;
assign v_19_out0 = A_366_out0[0:0];
assign v_75_out0 = A_366_out0[6:6];
assign v_99_out0 = A_366_out0[5:5];
assign v_125_out0 = A_366_out0[4:4];
assign v_165_out0 = A_366_out0[8:8];
assign v_215_out0 = A_366_out0[9:9];
assign v_294_out0 = A_366_out0[1:1];
assign v_299_out0 = A_366_out0[12:12];
assign v_318_out0 = A_366_out0[10:10];
assign v_331_out0 = A_366_out0[3:3];
assign v_383_out0 = A_366_out0[11:11];
assign v_485_out0 = A_366_out0[13:13];
assign XOR1_523_out0 = OP2_615_out0 ^ C1_544_out0;
assign v_581_out0 = A_366_out0[14:14];
assign v_596_out0 = A_366_out0[2:2];
assign v_616_out0 = A_366_out0[7:7];
assign v_638_out0 = A_366_out0[15:15];
assign G10_31_out0 = ! v_215_out0;
assign G13_116_out0 = ! v_299_out0;
assign G9_212_out0 = ! v_165_out0;
assign G12_216_out0 = ! v_383_out0;
assign G14_221_out0 = ! v_485_out0;
assign G5_253_out0 = ! v_125_out0;
assign G2_282_out0 = ! v_294_out0;
assign G16_314_out0 = ! v_638_out0;
assign G4_321_out0 = ! v_331_out0;
assign G15_351_out0 = ! v_581_out0;
assign G8_463_out0 = ! v_616_out0;
assign G7_536_out0 = ! v_75_out0;
assign G6_556_out0 = ! v_99_out0;
assign G3_582_out0 = ! v_596_out0;
assign MUX1_609_out0 = v_220_out0 ? XOR1_523_out0 : OP2_615_out0;
assign G11_619_out0 = ! v_318_out0;
assign G1_622_out0 = ! v_19_out0;
assign v_414_out0 = { G15_351_out0,G16_314_out0 };
assign {A1_597_out1,A1_597_out0 } = OP1_466_out0 + MUX1_609_out0 + MUX2_280_out0;
assign OUT_295_out0 = A1_597_out0;
assign v_317_out0 = { G14_221_out0,v_414_out0 };
assign v_329_out0 = A1_597_out0[15:15];
assign COUT_341_out0 = A1_597_out1;
assign CFF_11_out0 = v_329_out0;
assign MUX1_512_out0 = EQ1_535_out0 ? OP2_486_out0 : OUT_295_out0;
assign v_632_out0 = { G13_116_out0,v_317_out0 };
assign v_417_out0 = { G12_216_out0,v_632_out0 };
assign v_514_out0 = { G11_619_out0,v_417_out0 };
assign v_511_out0 = { G10_31_out0,v_514_out0 };
assign v_281_out0 = { G9_212_out0,v_511_out0 };
assign v_234_out0 = { G8_463_out0,v_281_out0 };
assign v_332_out0 = { G7_536_out0,v_234_out0 };
assign v_79_out0 = { G6_556_out0,v_332_out0 };
assign v_623_out0 = { G5_253_out0,v_79_out0 };
assign v_412_out0 = { G4_321_out0,v_623_out0 };
assign v_145_out0 = { G3_582_out0,v_412_out0 };
assign v_48_out0 = { G2_282_out0,v_145_out0 };
assign v_423_out0 = { G1_622_out0,v_48_out0 };
assign Y_12_out0 = v_423_out0;
assign MUX3_340_out0 = EQ5_277_out0 ? Y_12_out0 : OP2_486_out0;
assign B_464_out0 = MUX3_340_out0;
assign v_45_out0 = B_464_out0[1:1];
assign v_180_out0 = B_464_out0[15:15];
assign v_199_out0 = B_464_out0[2:2];
assign v_224_out0 = B_464_out0[11:11];
assign v_264_out0 = B_464_out0[9:9];
assign v_323_out0 = B_464_out0[14:14];
assign v_360_out0 = B_464_out0[13:13];
assign v_435_out0 = B_464_out0[10:10];
assign v_447_out0 = B_464_out0[5:5];
assign v_487_out0 = B_464_out0[12:12];
assign v_492_out0 = B_464_out0[8:8];
assign v_495_out0 = B_464_out0[6:6];
assign v_501_out0 = B_464_out0[4:4];
assign v_507_out0 = B_464_out0[3:3];
assign v_519_out0 = B_464_out0[7:7];
assign v_526_out0 = B_464_out0[0:0];
assign G13_15_out0 = v_574_out0 && v_487_out0;
assign G16_98_out0 = v_287_out0 && v_180_out0;
assign G11_184_out0 = v_286_out0 && v_435_out0;
assign G2_322_out0 = v_480_out0 && v_45_out0;
assign G8_328_out0 = v_239_out0 && v_519_out0;
assign G6_346_out0 = v_78_out0 && v_447_out0;
assign G4_371_out0 = v_227_out0 && v_507_out0;
assign G7_449_out0 = v_312_out0 && v_495_out0;
assign G12_468_out0 = v_114_out0 && v_224_out0;
assign G5_472_out0 = v_196_out0 && v_501_out0;
assign G3_506_out0 = v_33_out0 && v_199_out0;
assign G15_518_out0 = v_441_out0 && v_323_out0;
assign G14_540_out0 = v_27_out0 && v_360_out0;
assign G1_560_out0 = v_526_out0 && v_302_out0;
assign G9_578_out0 = v_135_out0 && v_492_out0;
assign G10_605_out0 = v_517_out0 && v_264_out0;
assign v_396_out0 = { G15_518_out0,G16_98_out0 };
assign v_603_out0 = { G14_540_out0,v_396_out0 };
assign v_278_out0 = { G13_15_out0,v_603_out0 };
assign v_34_out0 = { G12_468_out0,v_278_out0 };
assign v_539_out0 = { G11_184_out0,v_34_out0 };
assign v_397_out0 = { G10_605_out0,v_539_out0 };
assign v_219_out0 = { G9_578_out0,v_397_out0 };
assign v_122_out0 = { G8_328_out0,v_219_out0 };
assign v_426_out0 = { G7_449_out0,v_122_out0 };
assign v_58_out0 = { G6_346_out0,v_426_out0 };
assign v_285_out0 = { G5_472_out0,v_58_out0 };
assign v_319_out0 = { G4_371_out0,v_285_out0 };
assign v_566_out0 = { G3_506_out0,v_319_out0 };
assign v_151_out0 = { G2_322_out0,v_566_out0 };
assign v_334_out0 = { G1_560_out0,v_151_out0 };
assign Y_599_out0 = v_334_out0;
assign MUX2_460_out0 = G8_470_out0 ? Y_599_out0 : MUX1_512_out0;
assign MUX4_231_out0 = EQ6_382_out0 ? Y_12_out0 : MUX2_460_out0;
assign ALUOUT_401_out0 = MUX4_231_out0;
assign MUX4_3_out0 = G2_542_out0 ? ALUOUT_401_out0 : REGDIN_551_out0;
assign ALUOUT_240_out0 = ALUOUT_401_out0;
assign ALUOUT_554_out0 = ALUOUT_401_out0;
assign EQ1_446_out0 = ALUOUT_554_out0 == 16'h0;
assign DIN3_461_out0 = MUX4_3_out0;
assign ALUOUT_503_out0 = ALUOUT_240_out0;


endmodule
